this is not a genuine template ;-)
